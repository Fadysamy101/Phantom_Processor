library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Reg is

    generic(
        address_bits : integer := 3; 
        word_width   : integer := 8   
    );
	 
    port(
        clk          : in std_logic;
        rst          : in std_logic;
        we           : in std_logic;  -- Write Enable
        write_address   : in std_logic_vector(address_bits-1 downto 0);
        read_address1   : in std_logic_vector(address_bits-1 downto 0);
        read_address2   : in std_logic_vector(address_bits-1 downto 0);
        data_in      : in std_logic_vector(word_width-1 downto 0);
        data_out1    : out std_logic_vector(word_width-1 downto 0);
        data_out2    : out std_logic_vector(word_width-1 downto 0)
    );
	 
end entity Reg;



architecture behavioral of Reg is

    type reg_array is array ((2**address_bits)-1 downto 0) of std_logic_vector(word_width-1 downto 0);
    signal REGISTERS : reg_array;

begin

    process(clk, rst)
    begin
	 
        if rst = '1' then
            
            for i in 0 to (2**address_bits)-1 loop
				
                REGISTERS(i) <= (others => '0');
					 
            end loop;
				

        elsif rising_edge(clk) then
		  
            if we = '1' then
				
                REGISTERS(to_integer(unsigned(write_address))) <= data_in;
					 
            end if;
				
        end if;
    end process;
	 
	 

    data_out1 <= REGISTERS(to_integer(unsigned(read_address1)));
    data_out2 <= REGISTERS(to_integer(unsigned(read_address2)));

end architecture behavioral;
